RC or RL Lowpass Filter
*Lowpass Filter
*Student: Jose Lopez

vin 1 0 dc 0 ac 1      ;AC Source

*First circuit

*c1 2 0 200nf                ;Capacitance
*r1 1 2 1k                   ;Resistance

*Second circuit
r2 2 0 1000                     ;Resistance
l1 1 2 200mh                    ;Inductance

.control
*AC analysis from 1 Hz to 10 KHz
ac dec 1000 1 100k 
gnuplot Filter v(2)                     ;Plot gain
gnuplot Filter2 vdb(2)                  ;Plot gain in db
gnuplot Filter3 phase(v(2))             ;Plot phase  
.endc 
.end 