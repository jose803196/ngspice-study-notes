RC o RL Highpass Filter
*Highpass Filter
*Student: Jose Lopez

vin 1 0 dc 0 ac 1      ;AC Source

*First circuit

*c1 1 2 200nf                ;Capacitance
*r1 2 0 1k                   ;Resistance

*Second circuit
r2 1 2 1000                     ;Resistance
l1 2 0 200mh                    ;Inductance

.control
*AC analysis from 1 KHz to 10 KHz
ac dec 1000 1 100k 
gnuplot Filter v(2)                     ;Plot gain
gnuplot Filter2 vdb(2)                  ;Plot gain in db
gnuplot Filter3 phase(v(2))             ;Plot phase  
.endc 
.end 